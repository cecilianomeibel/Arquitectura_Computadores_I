module Adder(
    input logic [11:0]  a,b,
	 output logic [11:0] c
);

    assign c = a + b;

endmodule