module Adder(
    input logic [14:0]  a,b,
	 output logic [14:0] c
);

    assign c = a + b;

endmodule